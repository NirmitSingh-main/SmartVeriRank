module test;
initial begin
$display("Verilog working!");
$finish;
end
endmodule

